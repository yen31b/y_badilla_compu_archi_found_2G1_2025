module UART_top(
	 input  logic clk,
    input  logic rst,
    input  logic uart_rx,
    output logic uart_tx
);

	